
module niosii_top (
	clk_1_clk,
	reset_1_reset_n);	

	input		clk_1_clk;
	input		reset_1_reset_n;
endmodule
