
module niosii_top (
	clk_1_clk,
	pio_0_external_connection_export,
	reset_1_reset_n);	

	input		clk_1_clk;
	output	[9:0]	pio_0_external_connection_export;
	input		reset_1_reset_n;
endmodule
